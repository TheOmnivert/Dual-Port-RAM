///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Created by : Gourav Chandra Naidu
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
class dpram_sequence extends uvm_sequence

	function new(string name);
		super.new(name,this);
	endfunction
	
	task body();
		
	endtask
	
	
endclass