class dpram_driver extends uvm_driver
	
	`uvm_component_utils(dpram_driver)
	
	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction
	
	function void build_phase(phase);
	
	endfunction
	
endclass